module full_adder(
input a,
input b,
input cin,
output sum,
output cout);

module rca_4bit(a,b,c,s,carry);
input [3:0]a,b;
input c;
output [3:0]s;
output carry;





endmodule
